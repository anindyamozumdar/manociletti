`timescale 1ns/100ps

module Circuit_ex_03_31_a (A, B, C, D, F);

  output F;
  input A, B, C, D;
  wire w1, w2, w3, w4, w5;

  and G1 (w1, C, D);
  or G2 (w2, w1, B);
  and G3 (w3, w2, A);
  not G4 (w4, C);
  and G5 (w5, w4, B);
  or G6 (F, w3, w5);

endmodule
